module uart_top_tb(
    
);

    reg clk;
    reg rxd;
    reg txd;

endmodule